* Spice description of alu3b7_cougar
* Spice driver version -1217853383
* Date ( dd/mm/yyyy hh:mm:ss ): 22/04/2018 at 15:37:11

* INTERF a[0] a[1] a[2] b[0] b[1] b[2] resultado[0] resultado[1] 
* INTERF resultado[2] resultado[3] resultado[4] resultado[5] s[0] s[1] s[2] 
* INTERF vdd vss 


.subckt alu3b7_cougar 242 267 396 278 269 376 395 384 381 370 367 359 373 350 
+ 401 403 353 
* NET 13 = na2_x1_3_sig
* NET 18 = na3_x1_2_sig
* NET 20 = o2_x2_sig
* NET 22 = o2_x2_2_sig
* NET 36 = not_aux3
* NET 39 = inv_x2_3_sig
* NET 40 = not_aux32
* NET 42 = noa22_x1_2_sig
* NET 47 = a2_x2_7_sig
* NET 48 = o2_x2_3_sig
* NET 59 = inv_x2_7_sig
* NET 62 = not_aux17
* NET 65 = aux37
* NET 66 = a2_x2_5_sig
* NET 67 = no2_x1_3_sig
* NET 70 = aux33
* NET 72 = a3_x2_4_sig
* NET 81 = ao22_x2_sig
* NET 82 = a2_x2_4_sig
* NET 86 = no2_x1_2_sig
* NET 87 = not_aux14
* NET 95 = aux36
* NET 96 = no2_x1_6_sig
* NET 104 = an12_x1_sig
* NET 109 = oa2ao222_x2_sig
* NET 112 = oa2a22_x2_5_sig
* NET 113 = nao2o22_x1_2_sig
* NET 119 = no2_x1_4_sig
* NET 122 = ao22_x2_5_sig
* NET 123 = ao22_x2_4_sig
* NET 125 = a2_x2_6_sig
* NET 131 = not_aux23
* NET 134 = not_aux18
* NET 135 = no3_x1_4_sig
* NET 136 = oa2ao222_x2_2_sig
* NET 141 = not_aux33
* NET 149 = aux34
* NET 157 = a3_x2_sig
* NET 161 = a2_x2_sig
* NET 163 = a2_x2_2_sig
* NET 170 = a2_x2_3_sig
* NET 171 = not_aux4
* NET 175 = noa22_x1_sig
* NET 177 = not_aux6
* NET 179 = nao22_x1_sig
* NET 180 = not_a[0]
* NET 198 = inv_x2_4_sig
* NET 199 = not_aux35
* NET 202 = not_aux21
* NET 205 = not_aux7
* NET 211 = not_b[1]
* NET 212 = not_aux1
* NET 219 = not_aux0
* NET 220 = na3_x1_sig
* NET 225 = not_aux5
* NET 227 = na2_x1_sig
* NET 231 = oa2a22_x2_sig
* NET 233 = aux1
* NET 242 = a[0]
* NET 246 = aux9
* NET 249 = xr2_x1_5_sig
* NET 252 = xr2_x1_4_sig
* NET 255 = aux12
* NET 257 = inv_x2_5_sig
* NET 258 = not_s[0]
* NET 261 = na2_x1_2_sig
* NET 263 = aux2
* NET 266 = inv_x2_sig
* NET 267 = a[1]
* NET 269 = b[1]
* NET 271 = xr2_x1_2_sig
* NET 274 = nxr2_x1_sig
* NET 278 = b[0]
* NET 279 = not_b[0]
* NET 280 = no2_x1_sig
* NET 294 = noa22_x1_3_sig
* NET 295 = inv_x2_6_sig
* NET 296 = no3_x1_sig
* NET 299 = no3_x1_2_sig
* NET 303 = not_a[1]
* NET 304 = not_aux22
* NET 308 = na3_x1_3_sig
* NET 312 = not_b[2]
* NET 313 = no3_x1_3_sig
* NET 315 = na2_x1_4_sig
* NET 318 = nao2o22_x1_3_sig
* NET 319 = a3_x2_5_sig
* NET 322 = o3_x2_sig
* NET 323 = ao22_x2_3_sig
* NET 324 = ao22_x2_2_sig
* NET 330 = no2_x1_5_sig
* NET 331 = a3_x2_2_sig
* NET 332 = nao2o22_x1_sig
* NET 337 = oa22_x2_sig
* NET 341 = xr2_x1_sig
* NET 343 = oa2a22_x2_2_sig
* NET 350 = s[1]
* NET 353 = vss
* NET 354 = not_aux30
* NET 355 = aux38
* NET 356 = not_aux10
* NET 357 = o4_x2_sig
* NET 359 = resultado[5]
* NET 360 = a2_x2_8_sig
* NET 361 = inv_x2_8_sig
* NET 364 = na2_x1_5_sig
* NET 367 = resultado[4]
* NET 369 = aux31
* NET 370 = resultado[3]
* NET 371 = inv_x2_2_sig
* NET 373 = s[0]
* NET 374 = aux13
* NET 375 = not_a[2]
* NET 376 = b[2]
* NET 378 = a3_x2_3_sig
* NET 380 = mx3_x2_sig
* NET 381 = resultado[2]
* NET 384 = resultado[1]
* NET 385 = oa22_x2_2_sig
* NET 389 = not_s[1]
* NET 390 = oa2a22_x2_3_sig
* NET 395 = resultado[0]
* NET 396 = a[2]
* NET 398 = xr2_x1_3_sig
* NET 400 = oa2a22_x2_4_sig
* NET 401 = s[2]
* NET 403 = vdd
* NET 404 = not_s[2]
Mtr_00770 404 401 403 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00769 403 371 372 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00768 378 372 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00767 403 401 372 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00766 372 374 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00765 387 391 392 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00764 403 386 393 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00763 388 389 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00762 392 385 388 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00761 393 398 387 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00760 394 390 393 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00759 392 404 394 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00758 381 392 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00757 391 404 403 403 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00756 403 389 386 403 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00755 403 382 385 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00754 383 378 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00753 383 380 382 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00752 382 404 383 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00751 379 374 377 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00750 379 375 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00749 403 376 379 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00748 377 396 379 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00747 390 377 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00746 374 376 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00745 403 373 374 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00744 397 396 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00743 403 400 402 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00742 398 397 399 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00741 399 400 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00740 399 402 398 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00739 403 396 399 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00738 375 396 403 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00737 368 375 369 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00736 403 373 368 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00735 371 369 403 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00734 403 354 359 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00733 358 357 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00732 359 360 358 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00731 366 361 365 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00730 362 373 366 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00729 363 364 362 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00728 403 356 363 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00727 403 365 357 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00726 364 396 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00725 403 376 364 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00724 361 355 403 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00723 403 334 337 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00722 288 331 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00721 288 332 334 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00720 334 404 288 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00719 293 389 355 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00718 403 401 293 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00717 389 350 403 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00716 292 342 347 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00715 403 336 291 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00714 289 389 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00713 347 337 289 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00712 291 341 292 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00711 290 343 291 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00710 347 404 290 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00709 384 347 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00708 342 404 403 403 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00707 403 389 336 403 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00706 370 326 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00705 286 324 285 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00704 286 330 403 403 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00703 403 322 286 403 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00702 285 323 326 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00701 326 355 286 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00700 403 308 311 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00699 319 311 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00698 403 369 311 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00697 311 315 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00696 287 350 330 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00695 403 401 287 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00694 315 312 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00693 403 356 315 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00692 403 313 283 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00691 283 319 284 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00690 284 318 320 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00689 322 320 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00688 403 304 308 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00687 308 303 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00686 308 312 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00685 295 355 403 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00684 403 354 367 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00683 281 294 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00682 367 295 281 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00681 360 305 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00680 403 303 305 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00679 305 304 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00678 403 296 354 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00677 282 375 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00676 354 299 282 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00675 279 278 403 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00674 266 263 403 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00673 273 271 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00672 403 280 277 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00671 341 273 276 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00670 276 280 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00669 276 277 341 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00668 403 271 276 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00667 263 269 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00666 403 373 263 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00665 275 274 280 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00664 403 279 275 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00663 403 261 262 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00662 331 262 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00661 403 401 262 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00660 262 263 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00659 268 267 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00658 403 269 272 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00657 271 268 270 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00656 270 269 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00655 270 272 271 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00654 403 267 270 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00653 261 267 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00652 403 258 261 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00651 264 263 265 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00650 264 269 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00649 403 303 264 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00648 265 267 264 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00647 343 265 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00646 251 249 250 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00645 251 267 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00644 403 252 251 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00643 250 303 251 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00642 400 250 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00641 403 303 260 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00640 259 257 313 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00639 260 312 259 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00638 257 255 403 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00637 253 376 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00636 403 255 256 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00635 252 253 254 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00634 254 255 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00633 254 256 252 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00632 403 376 254 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00631 245 376 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00630 403 246 247 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00629 249 245 248 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00628 248 246 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00627 248 247 249 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00626 403 376 248 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00625 403 240 196 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00624 196 241 274 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00623 196 242 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00622 274 373 196 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00621 403 242 241 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00620 240 373 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00619 403 278 220 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00618 220 258 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00617 220 401 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00616 191 279 223 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00615 403 242 191 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00614 225 223 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00613 194 232 237 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00612 403 226 195 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00611 192 350 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00610 237 227 192 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00609 195 231 194 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00608 193 233 195 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00607 237 401 193 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00606 395 237 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00605 232 401 403 403 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00604 403 350 226 403 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00603 227 219 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00602 403 220 227 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00601 403 350 186 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00600 187 202 296 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00599 186 401 187 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00598 212 233 403 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00597 403 356 189 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00596 255 225 189 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00595 189 373 255 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00594 211 269 403 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00593 403 205 188 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00592 246 258 188 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00591 188 212 246 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00590 356 209 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00589 403 212 209 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00588 209 211 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00587 198 246 403 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00586 318 198 185 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00585 185 199 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00584 184 396 318 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00583 403 202 184 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00582 182 258 181 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00581 182 279 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00580 403 373 182 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00579 181 180 182 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00578 231 181 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00577 403 225 179 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00576 178 177 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00575 179 180 178 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00574 403 266 176 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00573 175 179 176 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00572 176 258 175 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00571 233 183 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00570 403 278 183 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00569 183 242 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00568 205 166 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00567 403 225 166 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00566 166 211 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00565 170 173 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00564 403 258 173 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00563 173 219 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00562 403 167 168 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00561 168 169 219 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00560 168 242 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00559 219 278 168 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00558 403 242 169 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00557 167 278 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00556 332 175 174 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00555 174 303 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00554 172 267 332 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00553 403 171 172 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00552 155 312 156 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00551 403 267 155 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00550 199 156 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00549 403 205 164 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00548 162 161 299 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00547 164 312 162 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00546 403 258 158 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00545 158 163 159 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00544 159 157 160 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00543 202 160 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00542 163 165 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00541 403 205 165 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00540 165 312 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00539 105 141 119 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00538 403 211 105 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00537 153 269 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00536 403 233 152 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00535 131 153 128 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00534 128 233 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00533 128 152 131 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00532 403 269 128 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00531 403 145 123 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00530 145 303 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00529 403 125 120 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00528 120 119 145 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00527 403 146 323 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00526 146 396 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00525 403 122 124 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00524 124 123 146 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00523 125 147 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00522 403 149 147 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00521 147 131 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00520 136 101 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00519 97 96 98 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00518 97 95 403 403 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00517 403 304 97 403 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00516 98 104 101 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00515 101 267 97 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00514 113 170 107 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00513 107 312 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00512 106 279 113 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00511 403 141 106 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00510 77 118 115 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00509 403 111 78 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00508 75 396 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00507 115 109 75 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00506 78 112 77 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00505 79 113 78 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00504 115 267 79 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00503 380 115 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00502 118 267 403 403 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00501 403 396 111 403 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00500 103 149 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00499 403 103 102 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00498 102 131 104 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00497 403 312 132 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00496 157 132 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00495 403 134 132 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00494 132 267 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00493 161 133 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00492 403 134 133 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00491 133 267 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00490 403 135 93 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00489 294 136 93 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00488 93 396 294 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00487 92 199 95 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00486 403 373 92 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00485 87 88 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00484 403 279 88 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00483 88 269 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00482 82 80 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00481 403 180 80 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00480 80 269 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00479 403 83 81 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00478 83 149 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00477 403 86 84 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00476 84 82 83 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00475 85 87 86 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00474 403 180 85 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00473 109 73 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00472 76 72 74 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00471 76 242 403 403 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00470 403 95 76 403 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00469 74 81 73 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00468 73 267 76 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00467 403 70 71 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00466 72 71 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00465 403 269 71 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00464 71 212 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00463 403 171 61 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00462 60 59 135 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00461 61 312 60 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00460 58 303 65 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00459 403 396 58 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00458 64 304 67 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00457 403 141 64 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00456 59 65 403 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00455 403 69 324 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00454 69 65 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00453 403 66 68 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00452 68 67 69 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00451 63 141 96 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00450 403 62 63 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00449 403 43 122 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00448 43 267 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00447 403 42 26 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00446 26 47 43 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00445 403 39 23 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00444 42 48 23 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00443 23 40 42 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00442 30 87 49 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00441 403 242 30 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00440 48 49 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00439 47 46 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00438 403 70 46 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00437 46 87 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00436 39 149 403 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00435 303 267 403 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00434 62 278 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00433 403 269 62 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00432 12 36 33 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00431 403 373 12 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00430 171 33 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00429 17 180 38 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00428 403 278 17 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00427 40 38 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00426 14 312 149 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00425 403 373 14 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00424 11 62 32 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00423 403 180 11 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00422 304 32 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00421 10 62 31 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00420 403 242 10 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00419 134 31 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00418 66 37 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00417 403 149 37 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00416 37 36 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00415 403 27 29 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00414 29 28 177 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00413 29 278 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00412 177 269 29 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00411 403 278 28 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00410 27 269 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00409 141 70 403 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00408 258 373 403 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00407 9 373 70 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00406 403 376 9 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00405 16 18 15 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00404 16 70 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00403 403 13 16 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00402 15 376 16 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00401 112 15 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00400 13 36 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00399 403 177 13 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00398 19 40 21 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00397 403 269 19 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00396 20 21 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00395 36 242 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00394 403 269 36 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00393 403 258 18 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00392 18 20 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00391 18 22 403 403 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00390 25 177 24 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00389 403 242 25 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00388 22 24 403 403 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00387 312 376 403 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00386 180 242 403 403 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00385 353 401 404 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00384 353 372 378 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00383 316 371 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00382 317 374 316 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00381 372 401 317 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00380 353 404 391 353 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00379 386 389 353 353 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00378 349 398 340 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00377 340 404 392 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00376 392 391 348 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00375 348 390 349 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00374 353 389 349 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00373 339 386 353 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00372 392 385 339 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00371 353 392 381 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00370 385 382 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00369 353 378 382 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00368 335 380 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00367 382 404 335 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00366 329 374 377 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00365 353 396 329 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00364 327 375 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00363 377 376 327 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00362 353 377 390 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00361 353 376 321 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00360 321 373 374 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00359 402 400 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00358 353 396 397 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00357 351 397 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00356 398 402 351 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00355 352 396 398 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00354 353 400 352 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00353 353 396 375 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00352 369 373 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00351 353 375 369 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00350 353 369 371 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00349 298 357 359 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00348 359 360 298 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00347 298 354 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00346 365 356 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00345 353 361 365 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00344 353 364 365 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00343 365 373 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00342 357 365 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00341 353 396 302 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00340 302 376 364 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00339 353 355 361 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00338 337 334 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00337 353 331 334 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00336 333 332 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00335 334 404 333 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00334 355 401 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00333 353 389 355 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00332 353 350 389 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00331 353 404 342 353 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00330 336 389 353 353 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00329 344 341 345 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00328 345 404 347 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00327 347 342 346 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00326 346 343 344 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00325 353 389 344 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00324 338 336 353 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00323 347 337 338 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00322 353 347 384 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00321 353 326 370 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00320 353 323 328 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00319 328 324 353 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00318 326 330 325 353 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00317 325 322 353 353 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00316 328 355 326 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00315 353 311 319 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00314 309 308 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00313 310 315 309 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00312 311 369 310 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00311 330 401 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00310 353 350 330 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00309 353 312 314 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00308 314 356 315 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00307 320 318 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00306 320 313 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00305 353 319 320 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00304 353 320 322 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00303 353 312 307 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00302 307 304 306 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00301 306 303 308 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00300 353 355 295 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00299 297 294 367 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00298 367 295 297 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00297 297 354 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00296 305 304 301 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00295 353 305 360 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00294 301 303 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00293 300 375 354 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00292 354 299 300 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00291 300 296 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00290 353 278 279 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00289 353 263 266 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00288 277 280 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00287 353 271 273 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00286 238 273 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00285 341 277 238 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00284 239 271 341 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00283 353 280 239 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00282 353 269 221 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00281 221 373 263 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00280 280 279 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00279 353 274 280 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00278 353 262 331 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00277 217 261 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00276 218 263 217 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00275 262 401 218 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00274 272 269 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00273 353 267 268 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00272 230 268 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00271 271 272 230 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00270 229 267 271 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00269 353 269 229 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00268 353 267 214 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00267 214 258 261 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00266 224 263 265 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00265 353 267 224 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00264 222 269 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00263 265 303 222 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00262 353 265 343 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00261 203 249 250 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00260 353 303 203 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00259 204 267 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00258 250 252 204 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00257 353 250 400 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00256 353 312 313 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00255 313 303 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00254 313 257 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00253 353 255 257 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00252 256 255 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00251 353 376 253 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00250 207 253 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00249 252 256 207 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00248 208 376 252 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00247 353 255 208 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00246 247 246 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00245 353 376 245 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00244 197 245 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00243 249 247 197 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00242 201 376 249 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00241 353 246 201 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00240 353 242 244 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00239 244 240 274 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00238 274 241 243 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00237 243 373 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00236 353 373 240 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00235 241 242 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00234 353 401 216 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00233 216 278 215 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00232 215 258 220 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00231 225 223 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00230 223 242 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00229 353 279 223 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00228 353 401 232 353 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00227 226 350 353 353 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00226 236 231 235 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00225 235 401 237 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00224 237 232 234 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00223 234 233 236 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00222 353 350 236 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00221 228 226 353 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00220 237 227 228 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00219 353 237 395 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00218 353 219 190 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00217 190 220 227 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00216 353 401 296 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00215 296 350 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00214 296 202 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00213 353 233 212 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00212 353 225 210 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00211 210 373 255 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00210 255 356 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00209 353 269 211 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00208 353 258 206 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00207 206 212 246 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00206 246 205 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00205 209 211 213 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00204 353 209 356 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00203 213 212 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00202 353 246 198 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00201 353 202 200 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00200 200 396 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00199 318 198 200 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00198 200 199 318 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00197 151 258 181 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00196 353 180 151 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00195 150 279 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00194 181 373 150 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00193 353 181 231 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00192 148 177 179 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00191 179 180 148 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00190 148 225 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00189 353 179 144 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00188 144 258 175 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00187 175 266 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00186 183 242 154 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00185 353 183 233 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00184 154 278 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00183 166 211 138 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00182 353 166 205 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00181 138 225 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00180 173 219 142 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00179 353 173 170 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00178 142 258 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00177 353 242 140 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00176 140 167 219 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00175 219 169 139 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00174 139 278 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00173 353 278 167 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00172 169 242 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00171 353 171 143 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00170 143 267 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00169 332 175 143 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00168 143 303 332 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00167 199 156 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00166 156 267 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00165 353 312 156 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00164 353 312 299 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00163 299 205 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00162 299 161 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00161 160 157 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00160 160 258 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00159 353 163 160 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00158 353 160 202 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00157 165 312 137 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00156 353 165 163 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00155 137 205 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00154 119 211 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00153 353 141 119 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00152 152 233 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00151 353 269 153 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00150 130 153 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00149 131 152 130 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00148 129 269 131 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00147 353 233 129 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00146 145 125 121 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00145 121 119 145 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00144 353 303 121 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00143 123 145 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00142 146 122 126 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00141 126 123 146 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00140 353 396 126 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00139 323 146 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00138 147 131 127 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00137 353 147 125 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00136 127 149 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00135 353 101 136 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00134 353 104 100 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00133 100 96 353 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00132 101 95 99 353 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00131 99 304 353 353 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00130 100 267 101 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00129 353 141 108 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00128 108 279 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00127 113 170 108 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00126 108 312 113 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00125 353 267 118 353 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00124 111 396 353 353 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00123 116 112 114 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00122 114 267 115 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00121 115 118 117 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00120 117 113 116 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00119 353 396 116 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00118 110 111 353 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00117 115 109 110 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00116 353 115 380 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00115 353 149 103 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00114 104 103 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00113 353 131 104 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00112 353 132 157 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00111 90 312 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00110 89 267 90 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00109 132 134 89 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00108 133 267 91 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00107 353 133 161 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00106 91 134 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00105 353 136 94 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00104 94 396 294 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00103 294 135 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00102 95 373 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00101 353 199 95 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00100 88 269 57 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00099 353 88 87 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00098 57 279 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00097 80 269 55 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00096 353 80 82 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00095 55 180 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00094 83 86 56 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00093 56 82 83 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00092 353 149 56 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00091 81 83 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00090 86 180 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00089 353 87 86 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00088 353 73 109 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00087 353 81 53 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00086 53 72 353 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00085 73 242 54 353 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00084 54 95 353 353 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00083 53 267 73 353 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00082 353 71 72 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00081 51 70 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00080 52 212 51 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00079 71 269 52 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00078 353 312 135 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00077 135 171 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00076 135 59 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00075 65 396 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00074 353 303 65 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00073 67 141 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00072 353 304 67 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00071 353 65 59 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00070 69 66 50 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00069 50 67 69 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00068 353 65 50 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00067 324 69 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00066 96 62 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00065 353 141 96 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00064 43 42 44 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00063 44 47 43 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00062 353 267 44 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00061 122 43 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00060 353 48 41 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00059 41 40 42 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00058 42 39 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00057 48 49 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00056 49 242 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00055 353 87 49 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00054 46 87 45 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00053 353 46 47 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00052 45 70 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00051 353 149 39 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00050 353 267 303 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00049 353 278 34 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00048 34 269 62 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00047 171 33 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00046 33 373 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00045 353 36 33 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00044 40 38 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00043 38 278 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00042 353 180 38 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00041 149 373 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00040 353 312 149 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00039 304 32 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00038 32 180 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00037 353 62 32 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00036 134 31 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00035 31 242 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00034 353 62 31 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00033 37 36 35 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00032 353 37 66 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00031 35 149 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00030 353 278 8 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00029 8 27 177 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00028 177 28 7 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00027 7 269 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00026 353 269 27 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00025 28 278 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00024 353 70 141 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00023 353 373 258 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00022 70 376 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00021 353 373 70 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00020 4 18 15 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00019 353 376 4 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00018 3 70 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00017 15 13 3 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00016 353 15 112 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00015 353 36 2 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00014 2 177 13 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00013 20 21 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00012 21 269 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00011 353 40 21 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00010 353 242 1 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00009 1 269 36 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00008 353 22 6 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00007 6 258 5 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00006 5 20 18 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00005 22 24 353 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00004 24 242 353 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00003 353 177 24 353 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00002 353 376 312 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00001 353 242 180 353 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
C399 13 353 5.361e-14
C397 15 353 2.445e-14
C396 16 353 7.43e-15
C394 18 353 5.175e-14
C392 20 353 5.156e-14
C391 21 353 1.8635e-14
C390 22 353 6.091e-14
C389 23 353 6.05e-15
C388 24 353 1.8635e-14
C385 27 353 2.596e-14
C384 28 353 2.16e-14
C383 29 353 7.76e-15
C380 31 353 1.8635e-14
C379 32 353 1.8635e-14
C378 33 353 1.8635e-14
C375 36 353 1.1427e-13
C374 37 353 1.8635e-14
C373 38 353 1.8635e-14
C372 39 353 5.319e-14
C371 40 353 9.21e-14
C369 42 353 5.227e-14
C368 43 353 1.853e-14
C367 44 353 4.11e-15
C365 46 353 1.8635e-14
C364 47 353 4.889e-14
C363 48 353 6.311e-14
C362 49 353 1.8635e-14
C361 50 353 4.11e-15
C358 53 353 4.11e-15
C355 56 353 4.11e-15
C351 59 353 5.874e-14
C348 62 353 1.211e-13
C345 65 353 1.0728e-13
C344 66 353 5.233e-14
C343 67 353 5.297e-14
C341 69 353 1.853e-14
C340 70 353 2.2716e-13
C339 71 353 2.605e-14
C338 72 353 5.19e-14
C337 73 353 2.299e-14
C334 76 353 8.58e-15
C332 78 353 7.56e-15
C330 80 353 1.8635e-14
C329 81 353 5.702e-14
C328 82 353 5.489e-14
C327 83 353 1.853e-14
C324 86 353 4.921e-14
C323 87 353 1.0702e-13
C322 88 353 1.8635e-14
C317 93 353 6.05e-15
C315 95 353 1.2653e-13
C314 96 353 4.846e-14
C313 97 353 8.58e-15
C310 100 353 4.11e-15
C309 101 353 2.299e-14
C307 103 353 1.677e-14
C306 104 353 4.828e-14
C302 108 353 7.43e-15
C301 109 353 5.93e-14
C299 111 353 2.378e-14
C298 112 353 9.224e-14
C297 113 353 5e-14
C295 115 353 3.608e-14
C294 116 353 7.56e-15
C292 118 353 2.128e-14
C291 119 353 7.457e-14
C289 121 353 4.11e-15
C288 122 353 6.917e-14
C287 123 353 5.733e-14
C285 125 353 4.993e-14
C284 126 353 4.11e-15
C281 128 353 9.7e-15
C278 131 353 1.3249e-13
C277 132 353 2.605e-14
C276 133 353 1.8635e-14
C275 134 353 9.416e-14
C274 135 353 5.719e-14
C273 136 353 4.179e-14
C268 141 353 1.68e-13
C266 143 353 7.43e-15
C264 145 353 1.853e-14
C263 146 353 1.853e-14
C262 147 353 1.8635e-14
C261 148 353 4.11e-15
C260 149 353 2.5651e-13
C257 152 353 2.16e-14
C256 153 353 2.596e-14
C252 156 353 1.8635e-14
C251 157 353 6.315e-14
C248 160 353 2.455e-14
C247 161 353 5.938e-14
C245 163 353 4.933e-14
C243 165 353 1.8635e-14
C242 166 353 1.8635e-14
C241 167 353 2.596e-14
C240 168 353 7.76e-15
C239 169 353 2.16e-14
C238 170 353 5.713e-14
C237 171 353 1.5315e-13
C235 173 353 1.8635e-14
C233 175 353 4.747e-14
C232 176 353 6.05e-15
C231 177 353 2.0046e-13
C229 179 353 4.547e-14
C228 180 353 3.0795e-13
C227 181 353 2.445e-14
C226 182 353 7.43e-15
C225 183 353 1.8635e-14
C220 188 353 6.05e-15
C219 189 353 6.05e-15
C213 195 353 7.56e-15
C211 196 353 7.76e-15
C209 198 353 4.929e-14
C208 199 353 1.0389e-13
C207 200 353 7.43e-15
C205 202 353 8.736e-14
C202 205 353 1.1901e-13
C198 209 353 1.8635e-14
C196 211 353 1.1736e-13
C195 212 353 1.7279e-13
C188 219 353 8.684e-14
C187 220 353 5.75e-14
C184 223 353 1.8635e-14
C182 225 353 1.6359e-13
C181 226 353 2.378e-14
C180 227 353 6.932e-14
C176 231 353 4.784e-14
C175 232 353 2.128e-14
C174 233 353 1.5148e-13
C171 236 353 7.56e-15
C170 237 353 3.608e-14
C167 240 353 2.596e-14
C166 241 353 2.16e-14
C165 242 353 5.0582e-13
C161 245 353 2.596e-14
C160 246 353 1.0662e-13
C159 247 353 2.16e-14
C158 248 353 9.7e-15
C157 249 353 5.485e-14
C156 250 353 2.445e-14
C155 251 353 7.43e-15
C154 252 353 5.365e-14
C153 253 353 2.596e-14
C152 254 353 9.7e-15
C151 255 353 8.814e-14
C150 256 353 2.16e-14
C149 257 353 4.914e-14
C148 258 353 4.21391e-13
C145 261 353 4.761e-14
C144 262 353 2.605e-14
C143 263 353 1.0513e-13
C142 264 353 7.43e-15
C141 265 353 2.445e-14
C140 266 353 6.639e-14
C139 267 353 5.9443e-13
C138 268 353 2.596e-14
C137 269 353 5.7134e-13
C136 270 353 9.7e-15
C135 271 353 5.995e-14
C134 272 353 2.16e-14
C133 273 353 2.596e-14
C132 274 353 5.574e-14
C130 276 353 9.7e-15
C129 277 353 2.16e-14
C128 278 353 4.2344e-13
C127 279 353 2.7769e-13
C126 280 353 5.577e-14
C120 286 353 8.58e-15
C118 288 353 6.05e-15
C115 291 353 7.56e-15
C111 294 353 9.733e-14
C110 295 353 4.809e-14
C109 296 353 7.567e-14
C108 297 353 4.11e-15
C107 298 353 4.11e-15
C106 299 353 8.257e-14
C105 300 353 4.11e-15
C102 303 353 3.9884e-13
C101 304 353 2.1941e-13
C100 305 353 1.8635e-14
C97 308 353 5.295e-14
C94 311 353 2.605e-14
C93 312 353 4.8008e-13
C92 313 353 5.797e-14
C90 315 353 4.551e-14
C87 318 353 1.0067e-13
C86 319 353 5.925e-14
C85 320 353 2.455e-14
C83 322 353 6.032e-14
C82 323 353 1.1342e-13
C81 324 353 1.145e-13
C79 326 353 2.299e-14
C77 328 353 4.11e-15
C75 330 353 4.561e-14
C74 331 353 8.141e-14
C73 332 353 8.657e-14
C71 334 353 1.767e-14
C69 336 353 2.378e-14
C68 337 353 5.998e-14
C64 341 353 5.246e-14
C63 342 353 2.128e-14
C62 343 353 7.336e-14
C61 344 353 7.56e-15
C58 347 353 3.608e-14
C56 349 353 7.56e-15
C55 350 353 3.2669e-13
C52 353 353 4.61908e-12
C51 354 353 8.966e-14
C50 355 353 2.1574e-13
C49 356 353 1.636e-13
C48 357 353 4.459e-14
C46 359 353 3.04e-14
C45 360 353 6.121e-14
C44 361 353 5.619e-14
C41 364 353 4.821e-14
C40 365 353 2.72e-14
C38 367 353 6.232e-14
C36 369 353 7.942e-14
C35 370 353 4.664e-14
C34 371 353 4.959e-14
C33 372 353 2.605e-14
C32 373 353 6.5862e-13
C31 374 353 8.382e-14
C30 375 353 1.4234e-13
C29 376 353 4.7094e-13
C28 377 353 2.445e-14
C27 378 353 7.781e-14
C26 379 353 7.43e-15
C25 380 353 1.1019e-13
C24 381 353 4.202e-14
C23 382 353 1.767e-14
C22 383 353 6.05e-15
C21 384 353 4.226e-14
C20 385 353 6.118e-14
C19 386 353 2.378e-14
C16 389 353 1.406e-13
C15 390 353 7.336e-14
C14 391 353 2.128e-14
C13 392 353 3.608e-14
C12 393 353 7.56e-15
C10 395 353 8.306e-14
C9 396 353 5.6937e-13
C8 397 353 2.596e-14
C7 398 353 5.006e-14
C6 399 353 9.7e-15
C5 400 353 1.5753e-13
C4 401 353 3.8086e-13
C3 402 353 2.16e-14
C2 403 353 4.76805e-12
C1 404 353 1.757e-13
.ends alu3b7_cougar

